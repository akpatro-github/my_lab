magic
tech scmos
timestamp 1616527254
<< pwell >>
rect -26 -43 139 -6
<< nwell >>
rect -26 -6 139 31
<< polysilicon >>
rect -22 18 114 20
rect -22 8 -20 18
rect -15 13 22 15
rect -15 8 -13 13
rect -4 9 -2 11
rect 12 9 14 11
rect 20 9 22 13
rect 28 9 30 18
rect 80 14 110 16
rect 36 9 38 11
rect 40 9 42 11
rect 56 9 58 11
rect 72 9 74 11
rect 80 9 82 14
rect 88 10 106 12
rect 88 9 90 10
rect 104 9 106 10
rect 108 9 110 14
rect 112 9 114 18
rect 128 9 130 11
rect -4 -16 -2 3
rect 12 -16 14 3
rect 20 -16 22 3
rect 28 -16 30 3
rect 36 -16 38 3
rect 40 -16 42 3
rect 56 -4 58 3
rect 57 -8 58 -4
rect 56 -16 58 -8
rect 72 -16 74 3
rect 80 -16 82 3
rect 88 -16 90 3
rect 104 -16 106 3
rect 108 -16 110 3
rect 112 -16 114 3
rect 128 -4 130 3
rect 129 -8 130 -4
rect 128 -16 130 -8
rect -14 -30 -12 -21
rect -4 -24 -2 -22
rect 12 -30 14 -22
rect 20 -26 22 -22
rect 28 -24 30 -22
rect 36 -26 38 -22
rect 20 -28 38 -26
rect 40 -30 42 -22
rect 56 -24 58 -22
rect 72 -26 74 -22
rect 80 -24 82 -22
rect 88 -24 90 -22
rect 104 -26 106 -22
rect 72 -28 106 -26
rect 108 -30 110 -22
rect 112 -24 114 -22
rect 128 -24 130 -22
rect -14 -32 110 -30
<< ndiffusion >>
rect -9 -17 -4 -16
rect -5 -21 -4 -17
rect -9 -22 -4 -21
rect -2 -17 3 -16
rect -2 -21 -1 -17
rect -2 -22 3 -21
rect 7 -17 12 -16
rect 11 -21 12 -17
rect 7 -22 12 -21
rect 14 -17 20 -16
rect 14 -21 15 -17
rect 19 -21 20 -17
rect 14 -22 20 -21
rect 22 -17 28 -16
rect 22 -21 23 -17
rect 27 -21 28 -17
rect 22 -22 28 -21
rect 30 -17 36 -16
rect 30 -21 31 -17
rect 35 -21 36 -17
rect 30 -22 36 -21
rect 38 -22 40 -16
rect 42 -17 47 -16
rect 42 -21 43 -17
rect 42 -22 47 -21
rect 51 -17 56 -16
rect 55 -21 56 -17
rect 51 -22 56 -21
rect 58 -17 63 -16
rect 58 -21 59 -17
rect 58 -22 63 -21
rect 67 -17 72 -16
rect 71 -21 72 -17
rect 67 -22 72 -21
rect 74 -17 80 -16
rect 74 -21 75 -17
rect 79 -21 80 -17
rect 74 -22 80 -21
rect 82 -17 88 -16
rect 82 -21 83 -17
rect 87 -21 88 -17
rect 82 -22 88 -21
rect 90 -17 95 -16
rect 90 -21 91 -17
rect 90 -22 95 -21
rect 99 -17 104 -16
rect 103 -21 104 -17
rect 99 -22 104 -21
rect 106 -22 108 -16
rect 110 -22 112 -16
rect 114 -17 119 -16
rect 114 -21 115 -17
rect 114 -22 119 -21
rect 123 -17 128 -16
rect 127 -21 128 -17
rect 123 -22 128 -21
rect 130 -17 135 -16
rect 130 -21 131 -17
rect 130 -22 135 -21
<< pdiffusion >>
rect -9 8 -4 9
rect -5 4 -4 8
rect -9 3 -4 4
rect -2 8 3 9
rect -2 4 -1 8
rect -2 3 3 4
rect 7 8 12 9
rect 11 4 12 8
rect 7 3 12 4
rect 14 8 20 9
rect 14 4 15 8
rect 19 4 20 8
rect 14 3 20 4
rect 22 8 28 9
rect 22 4 23 8
rect 27 4 28 8
rect 22 3 28 4
rect 30 8 36 9
rect 30 4 31 8
rect 35 4 36 8
rect 30 3 36 4
rect 38 3 40 9
rect 42 8 47 9
rect 42 4 43 8
rect 42 3 47 4
rect 51 8 56 9
rect 55 4 56 8
rect 51 3 56 4
rect 58 8 63 9
rect 58 4 59 8
rect 58 3 63 4
rect 67 8 72 9
rect 71 4 72 8
rect 67 3 72 4
rect 74 8 80 9
rect 74 4 75 8
rect 79 4 80 8
rect 74 3 80 4
rect 82 8 88 9
rect 82 4 83 8
rect 87 4 88 8
rect 82 3 88 4
rect 90 8 95 9
rect 90 4 91 8
rect 90 3 95 4
rect 99 8 104 9
rect 103 4 104 8
rect 99 3 104 4
rect 106 3 108 9
rect 110 3 112 9
rect 114 8 119 9
rect 114 4 115 8
rect 114 3 119 4
rect 123 8 128 9
rect 127 4 128 8
rect 123 3 128 4
rect 130 8 135 9
rect 130 4 131 8
rect 130 3 135 4
<< metal1 >>
rect -26 24 7 28
rect 11 24 139 28
rect 7 15 10 24
rect 83 15 86 24
rect 0 12 18 15
rect 0 8 3 12
rect 15 8 18 12
rect 24 12 47 15
rect 24 8 27 12
rect 44 8 47 12
rect -26 4 -23 8
rect -16 1 -12 4
rect -26 -3 -12 1
rect 51 12 70 15
rect 51 8 54 12
rect 67 8 70 12
rect 75 12 95 15
rect 75 8 78 12
rect 92 8 95 12
rect 123 8 126 24
rect -9 -6 -6 4
rect 7 1 10 4
rect 24 1 27 4
rect 7 -2 27 1
rect -26 -10 -6 -6
rect 32 -5 35 4
rect 2 -8 53 -5
rect 60 -5 63 4
rect 67 1 70 4
rect 84 1 87 4
rect 99 1 102 4
rect 67 -2 102 1
rect 116 -5 119 4
rect 132 -4 135 4
rect 60 -8 125 -5
rect 132 -8 139 -4
rect -9 -17 -6 -10
rect 7 -14 27 -11
rect 7 -17 10 -14
rect 24 -17 27 -14
rect 32 -17 35 -8
rect 60 -17 63 -8
rect 116 -11 119 -8
rect 68 -14 87 -11
rect 68 -17 71 -14
rect 84 -17 87 -14
rect 99 -14 119 -11
rect 99 -17 102 -14
rect 132 -17 135 -8
rect -20 -21 -16 -17
rect 0 -36 3 -21
rect 16 -36 19 -21
rect 44 -36 47 -21
rect 51 -24 54 -21
rect 68 -24 71 -21
rect 51 -27 71 -24
rect 76 -36 79 -21
rect 92 -36 95 -21
rect 116 -24 119 -21
rect 123 -24 126 -21
rect 116 -27 126 -24
rect -26 -40 7 -36
rect 11 -40 139 -36
<< ntransistor >>
rect -4 -22 -2 -16
rect 12 -22 14 -16
rect 20 -22 22 -16
rect 28 -22 30 -16
rect 36 -22 38 -16
rect 40 -22 42 -16
rect 56 -22 58 -16
rect 72 -22 74 -16
rect 80 -22 82 -16
rect 88 -22 90 -16
rect 104 -22 106 -16
rect 108 -22 110 -16
rect 112 -22 114 -16
rect 128 -22 130 -16
<< ptransistor >>
rect -4 3 -2 9
rect 12 3 14 9
rect 20 3 22 9
rect 28 3 30 9
rect 36 3 38 9
rect 40 3 42 9
rect 56 3 58 9
rect 72 3 74 9
rect 80 3 82 9
rect 88 3 90 9
rect 104 3 106 9
rect 108 3 110 9
rect 112 3 114 9
rect 128 3 130 9
<< polycontact >>
rect -23 4 -19 8
rect -16 4 -12 8
rect -2 -8 2 -4
rect 53 -8 57 -4
rect 125 -8 129 -4
rect -16 -21 -12 -17
<< ndcontact >>
rect -9 -21 -5 -17
rect -1 -21 3 -17
rect 7 -21 11 -17
rect 15 -21 19 -17
rect 23 -21 27 -17
rect 31 -21 35 -17
rect 43 -21 47 -17
rect 51 -21 55 -17
rect 59 -21 63 -17
rect 67 -21 71 -17
rect 75 -21 79 -17
rect 83 -21 87 -17
rect 91 -21 95 -17
rect 99 -21 103 -17
rect 115 -21 119 -17
rect 123 -21 127 -17
rect 131 -21 135 -17
<< pdcontact >>
rect -9 4 -5 8
rect -1 4 3 8
rect 7 4 11 8
rect 15 4 19 8
rect 23 4 27 8
rect 31 4 35 8
rect 43 4 47 8
rect 51 4 55 8
rect 59 4 63 8
rect 67 4 71 8
rect 75 4 79 8
rect 83 4 87 8
rect 91 4 95 8
rect 99 4 103 8
rect 115 4 119 8
rect 123 4 127 8
rect 131 4 135 8
<< psubstratepcontact >>
rect 7 -40 11 -36
<< nsubstratencontact >>
rect 7 24 11 28
<< labels >>
rlabel metal1 -21 26 -21 26 4 VDD
rlabel metal1 -18 -38 -18 -38 1 GND
rlabel metal1 -18 -19 -18 -19 1 Cin
rlabel metal1 -23 -8 -23 -8 3 Cout
rlabel metal1 -22 -1 -22 -1 3 Bin
rlabel metal1 -25 6 -25 6 3 Ain
rlabel metal1 137 -6 137 -6 7 SUM
<< end >>
