* SPICE3 file created from /home/vlsi/Desktop/my_lab_logic/nand.ext - technology: scmos

.option scale=0.2u

M1000 GND B a_0_n21# GND nfet w=6 l=2
+  ad=30 pd=22 as=36 ps=24
M1001 VDD B out VDD pfet w=12 l=2
+  ad=120 pd=68 as=72 ps=36
M1002 a_0_n21# A out GND nfet w=6 l=2
+  ad=0 pd=0 as=30 ps=22
M1003 out A VDD VDD pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
C0 VDD GND 2.67fF
