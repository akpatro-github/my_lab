magic
tech scmos
timestamp 1602393362
<< nwell >>
rect -13 -8 22 24
<< ntransistor >>
rect -2 -21 0 -15
rect 6 -21 8 -15
<< ptransistor >>
rect -2 -2 0 10
rect 6 -2 8 10
<< ndiffusion >>
rect -7 -16 -2 -15
rect -3 -20 -2 -16
rect -7 -21 -2 -20
rect 0 -21 6 -15
rect 8 -17 13 -15
rect 8 -21 9 -17
<< pdiffusion >>
rect -7 6 -2 10
rect -3 2 -2 6
rect -7 -2 -2 2
rect 0 4 6 10
rect 0 0 1 4
rect 5 0 6 4
rect 0 -2 6 0
rect 8 6 13 10
rect 8 2 9 6
rect 8 -2 13 2
<< ndcontact >>
rect -7 -20 -3 -16
rect 9 -21 13 -17
<< pdcontact >>
rect -7 2 -3 6
rect 1 0 5 4
rect 9 2 13 6
<< psubstratepcontact >>
rect -9 -30 -5 -26
rect 1 -30 5 -26
rect 14 -30 18 -26
<< nsubstratencontact >>
rect -7 17 -3 21
rect 1 17 5 21
rect 9 17 13 21
<< polysilicon >>
rect -2 10 0 12
rect 6 10 8 12
rect -2 -10 0 -2
rect -10 -14 0 -10
rect -2 -15 0 -14
rect 6 -10 8 -2
rect 6 -14 9 -10
rect 6 -15 8 -14
rect -2 -23 0 -21
rect 6 -23 8 -21
<< polycontact >>
rect -14 -14 -10 -10
rect 9 -14 13 -10
<< metal1 >>
rect -13 17 -7 21
rect -3 17 1 21
rect 5 17 9 21
rect 13 17 22 21
rect -13 16 22 17
rect -7 6 -3 16
rect 9 6 13 16
rect 1 -9 5 0
rect -16 -14 -14 -10
rect -7 -13 5 -9
rect -7 -16 -3 -13
rect 13 -14 15 -10
rect 9 -26 13 -21
rect -12 -30 -9 -26
rect -5 -30 1 -26
rect 5 -30 14 -26
rect 18 -30 21 -26
rect -12 -31 21 -30
<< labels >>
rlabel psubstratepcontact 3 -28 3 -28 1 GND
rlabel nsubstratencontact 3 19 3 19 5 VDD
rlabel polycontact -12 -12 -12 -12 3 A
rlabel polycontact 11 -12 11 -12 1 B
rlabel metal1 3 -11 3 -11 1 out
<< end >>
